----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    03:27:31 10/21/2025 
-- Design Name: 
-- Module Name:    CIRCUITOSVhdlCircuito3_HSF - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity CIRCUITOSVhdlCircuito3_HSF is
    Port ( a : in  STD_LOGIC;
           b : in  STD_LOGIC;
           c : in  STD_LOGIC;
           d : in  STD_LOGIC;
			  negative_a : inout  STD_LOGIC;
			  negative_c : inout  STD_LOGIC;
			  t1 : inout  STD_LOGIC;
			  t2 : inout  STD_LOGIC;
			  t3 : inout  STD_LOGIC;
			  t4 : inout  STD_LOGIC;
			  t5 : inout  STD_LOGIC;
			  t6 : inout  STD_LOGIC;
			  t7 : inout  STD_LOGIC;
           s : out  STD_LOGIC);
end CIRCUITOSVhdlCircuito3_HSF;

architecture Behavioral of CIRCUITOSVhdlCircuito3_HSF is

begin
--Entries variations
negative_a<=not a;
negative_c<=not c;

--First column
t1<=b or d;
t2<=a and negative_c and d;
t3<=negative_a or b or negative_c;

--Second column
t4<=(not t2) or (not t3);

--Third column
t5<=c and (not t4);
t6<=(not t3) and d;

--Final
t7<=t1 or t5 or (not t6);
s<=not t7;

end Behavioral;

